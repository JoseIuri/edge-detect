`ifndef STOCHASTIC_TYPES
`define STOCHASTIC_TYPES

`endif